library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.perceptron_utility_pkg.all;

entity SigmoidLUT is
	port(
		x : IN std_logic_vector(BitO-1 downto 0);
		y : OUT std_logic_vector(BitY-1 downto 0);
		-- Basic Pins
		clk : IN std_logic;
		resetn : IN std_logic
	);

end SigmoidLUT;

architecture internal of SigmoidLUT is

	type SigmoidLUT_T is array(natural range<>) of natural;
	
	constant SigmoidLUT : SigmoidLUT_T :=(0, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 328, 329, 330, 331, 332, 333, 334, 335, 336, 336, 337, 338, 339, 340, 341, 342, 343, 344, 344, 345, 346, 347, 348, 349, 350, 351, 352, 352, 353, 354, 355, 356, 357, 358, 359, 359, 360, 361, 362, 363, 364, 365, 366, 366, 367, 368, 369, 370, 371, 372, 373, 373, 374, 375, 376, 377, 378, 379, 379, 380, 381, 382, 383, 384, 385, 385, 386, 387, 388, 389, 390, 391, 391, 392, 393, 394, 395, 396, 397, 397, 398, 399, 400, 401, 402, 403, 403, 404, 405, 406, 407, 408, 408, 409, 410, 411, 412, 413, 413, 414, 415, 416, 417, 418, 418, 419, 420, 421, 422, 423, 423, 424, 425, 426, 427, 428, 428, 429, 430, 431, 432, 433, 433, 434, 435, 436, 437, 437, 438, 439, 440, 441, 442, 442, 443, 444, 445, 446, 446, 447, 448, 449, 450, 450, 451, 452, 453, 454, 454, 455, 456, 457, 458, 458, 459, 460, 461, 462, 462, 463, 464, 465, 466, 466, 467, 468, 469, 470, 470, 471, 472, 473, 473, 474, 475, 476, 477, 477, 478, 479, 480, 481, 481, 482, 483, 484, 484, 485, 486, 487, 488, 488, 489, 490, 491, 491, 492, 493, 494, 494, 495, 496, 497, 498, 498, 499, 500, 501, 501, 502, 503, 504, 504, 505, 506, 507, 507, 508, 509, 510, 510, 511, 512, 513, 513, 514, 515, 516, 516, 517, 518, 519, 519, 520, 521, 522, 522, 523, 524, 525, 525, 526, 527, 527, 528, 529, 530, 530, 531, 532, 533, 533, 534, 535, 535, 536, 537, 538, 538, 539, 540, 541, 541, 542, 543, 543, 544, 545, 546, 546, 547, 548, 548, 549, 550, 551, 551, 552, 553, 553, 554, 555, 556, 556, 557, 558, 558, 559, 560, 560, 561, 562, 563, 563, 564, 565, 565, 566, 567, 567, 568, 569, 569, 570, 571, 572, 572, 573, 574, 574, 575, 576, 576, 577, 578, 578, 579, 580, 580, 581, 582, 582, 583, 584, 584, 585, 586, 587, 587, 588, 589, 589, 590, 591, 591, 592, 593, 593, 594, 595, 595, 596, 596, 597, 598, 598, 599, 600, 600, 601, 602, 602, 603, 604, 604, 605, 606, 606, 607, 608, 608, 609, 610, 610, 611, 611, 612, 613, 613, 614, 615, 615, 616, 617, 617, 618, 618, 619, 620, 620, 621, 622, 622, 623, 624, 624, 625, 625, 626, 627, 627, 628, 629, 629, 630, 630, 631, 632, 632, 633, 634, 634, 635, 635, 636, 637, 637, 638, 638, 639, 640, 640, 641, 641, 642, 643, 643, 644, 644, 645, 646, 646, 647, 648, 648, 649, 649, 650, 650, 651, 652, 652, 653, 653, 654, 655, 655, 656, 656, 657, 658, 658, 659, 659, 660, 661, 661, 662, 662, 663, 663, 664, 665, 665, 666, 666, 667, 667, 668, 669, 669, 670, 670, 671, 671, 672, 673, 673, 674, 674, 675, 675, 676, 677, 677, 678, 678, 679, 679, 680, 680, 681, 682, 682, 683, 683, 684, 684, 685, 685, 686, 687, 687, 688, 688, 689, 689, 690, 690, 691, 691, 692, 693, 693, 694, 694, 695, 695, 696, 696, 697, 697, 698, 698, 699, 700, 700, 701, 701, 702, 702, 703, 703, 704, 704, 705, 705, 706, 706, 707, 707, 708, 709, 709, 710, 710, 711, 711, 712, 712, 713, 713, 714, 714, 715, 715, 716, 716, 717, 717, 718, 718, 719, 719, 720, 720, 721, 721, 722, 722, 723, 723, 724, 724, 725, 725, 726, 726, 727, 727, 728, 728, 729, 729, 730, 730, 731, 731, 732, 732, 733, 733, 734, 734, 735, 735, 736, 736, 737, 737, 738, 738, 738, 739, 739, 740, 740, 741, 741, 742, 742, 743, 743, 744, 744, 745, 745, 746, 746, 747, 747, 747, 748, 748, 749, 749, 750, 750, 751, 751, 752, 752, 753, 753, 753, 754, 754, 755, 755, 756, 756, 757, 757, 758, 758, 758, 759, 759, 760, 760, 761, 761, 762, 762, 763, 763, 763, 764, 764, 765, 765, 766, 766, 766, 767, 767, 768, 768, 769, 769, 770, 770, 770, 771, 771, 772, 772, 773, 773, 773, 774, 774, 775, 775, 776, 776, 776, 777, 777, 778, 778, 779, 779, 779, 780, 780, 781, 781, 781, 782, 782, 783, 783, 784, 784, 784, 785, 785, 786, 786, 786, 787, 787, 788, 788, 788, 789, 789, 790, 790, 790, 791, 791, 792, 792, 792, 793, 793, 794, 794, 794, 795, 795, 796, 796, 796, 797, 797, 798, 798, 798, 799, 799, 800, 800, 800, 801, 801, 802, 802, 802, 803, 803, 803, 804, 804, 805, 805, 805, 806, 806, 807, 807, 807, 808, 808, 808, 809, 809, 810, 810, 810, 811, 811, 811, 812, 812, 813, 813, 813, 814, 814, 814, 815, 815, 815, 816, 816, 817, 817, 817, 818, 818, 818, 819, 819, 819, 820, 820, 821, 821, 821, 822, 822, 822, 823, 823, 823, 824, 824, 824, 825, 825, 825, 826, 826, 826, 827, 827, 828, 828, 828, 829, 829, 829, 830, 830, 830, 831, 831, 831, 832, 832, 832, 833, 833, 833, 834, 834, 834, 835, 835, 835, 836, 836, 836, 837, 837, 837, 838, 838, 838, 839, 839, 839, 840, 840, 840, 841, 841, 841, 842, 842, 842, 843, 843, 843, 844, 844, 844, 844, 845, 845, 845, 846, 846, 846, 847, 847, 847, 848, 848, 848, 849, 849, 849, 850, 850, 850, 850, 851, 851, 851, 852, 852, 852, 853, 853, 853, 854, 854, 854, 854, 855, 855, 855, 856, 856, 856, 857, 857, 857, 857, 858, 858, 858, 859, 859, 859, 860, 860, 860, 860, 861, 861, 861, 862, 862, 862, 862, 863, 863, 863, 864, 864, 864, 864, 865, 865, 865, 866, 866, 866, 866, 867, 867, 867, 868, 868, 868, 868, 869, 869, 869, 870, 870, 870, 870, 871, 871, 871, 871, 872, 872, 872, 873, 873, 873, 873, 874, 874, 874, 874, 875, 875, 875, 876, 876, 876, 876, 877, 877, 877, 877, 878, 878, 878, 878, 879, 879, 879, 880, 880, 880, 880, 881, 881, 881, 881, 882, 882, 882, 882, 883, 883, 883, 883, 884, 884, 884, 884, 885, 885, 885, 885, 886, 886, 886, 886, 887, 887, 887, 887, 888, 888, 888, 888, 889, 889, 889, 889, 890, 890, 890, 890, 891, 891, 891, 891, 892, 892, 892, 892, 893, 893, 893, 893, 893, 894, 894, 894, 894, 895, 895, 895, 895, 896, 896, 896, 896, 897, 897, 897, 897, 897, 898, 898, 898, 898, 899, 899, 899, 899, 900, 900, 900, 900, 900, 901, 901, 901, 901, 902, 902, 902, 902, 902, 903, 903, 903, 903, 904, 904, 904, 904, 904, 905, 905, 905, 905, 906, 906, 906, 906, 906, 907, 907, 907, 907, 907, 908, 908, 908, 908, 909, 909, 909, 909, 909, 910, 910, 910, 910, 910, 911, 911, 911, 911, 911, 912, 912, 912, 912, 913, 913, 913, 913, 913, 914, 914, 914, 914, 914, 915, 915, 915, 915, 915, 916, 916, 916, 916, 916, 917, 917, 917, 917, 917, 918, 918, 918, 918, 918, 918, 919, 919, 919, 919, 919, 920, 920, 920, 920, 920, 921, 921, 921, 921, 921, 922, 922, 922, 922, 922, 923, 923, 923, 923, 923, 923, 924, 924, 924, 924, 924, 925, 925, 925, 925, 925, 925, 926, 926, 926, 926, 926, 927, 927, 927, 927, 927, 927, 928, 928, 928, 928, 928, 929, 929, 929, 929, 929, 929, 930, 930, 930, 930, 930, 930, 931, 931, 931, 931, 931, 931, 932, 932, 932, 932, 932, 933, 933, 933, 933, 933, 933, 934, 934, 934, 934, 934, 934, 935, 935, 935, 935, 935, 935, 936, 936, 936, 936, 936, 936, 936, 937, 937, 937, 937, 937, 937, 938, 938, 938, 938, 938, 938, 939, 939, 939, 939, 939, 939, 940, 940, 940, 940, 940, 940, 940, 941, 941, 941, 941, 941, 941, 942, 942, 942, 942, 942, 942, 942, 943, 943, 943, 943, 943, 943, 944, 944, 944, 944, 944, 944, 944, 945, 945, 945, 945, 945, 945, 945, 946, 946, 946, 946, 946, 946, 946, 947, 947, 947, 947, 947, 947, 947, 948, 948, 948, 948, 948, 948, 948, 949, 949, 949, 949, 949, 949, 949, 950, 950, 950, 950, 950, 950, 950, 951, 951, 951, 951, 951, 951, 951, 952, 952, 952, 952, 952, 952, 952, 952, 953, 953, 953, 953, 953, 953, 953, 954, 954, 954, 954, 954, 954, 954, 954, 955, 955, 955, 955, 955, 955, 955, 955, 956, 956, 956, 956, 956, 956, 956, 957, 957, 957, 957, 957, 957, 957, 957, 958, 958, 958, 958, 958, 958, 958, 958, 958, 959, 959, 959, 959, 959, 959, 959, 959, 960, 960, 960, 960, 960, 960, 960, 960, 961, 961, 961, 961, 961, 961, 961, 961, 962, 962, 962, 962, 962, 962, 962, 962, 962, 963, 963, 963, 963, 963, 963, 963, 963, 963, 964, 964, 964, 964, 964, 964, 964, 964, 964, 965, 965, 965, 965, 965, 965, 965, 965, 965, 966, 966, 966, 966, 966, 966, 966, 966, 966, 967, 967, 967, 967, 967, 967, 967, 967, 967, 968, 968, 968, 968, 968, 968, 968, 968, 968, 968, 969, 969, 969, 969, 969, 969, 969, 969, 969, 970, 970, 970, 970, 970, 970, 970, 970, 970, 970, 971, 971, 971, 971, 971, 971, 971, 971, 971, 971, 972, 972, 972, 972, 972, 972, 972, 972, 972, 972, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 973, 974, 974, 974, 974, 974, 974, 974, 974, 974, 974, 975, 975, 975, 975, 975, 975, 975, 975, 975, 975, 975, 976, 976, 976, 976, 976, 976, 976, 976, 976, 976, 976, 977, 977, 977, 977, 977, 977, 977, 977, 977, 977, 977, 978, 978, 978, 978, 978, 978, 978, 978, 978, 978, 978, 978, 979, 979, 979, 979, 979, 979, 979, 979, 979, 979, 979, 979, 980, 980, 980, 980, 980, 980, 980, 980, 980, 980, 980, 980, 981, 981, 981, 981, 981, 981, 981, 981, 981, 981, 981, 981, 982, 982, 982, 982, 982, 982, 982, 982, 982, 982, 982, 982, 982, 983, 983, 983, 983, 983, 983, 983, 983, 983, 983, 983, 983, 984, 984, 984, 984, 984, 984, 984, 984, 984, 984, 984, 984, 984, 984, 985, 985, 985, 985, 985, 985, 985, 985, 985, 985, 985, 985, 985, 986, 986, 986, 986, 986, 986, 986, 986, 986, 986, 986, 986, 986, 986, 987, 987, 987, 987, 987, 987, 987, 987, 987, 987, 987, 987, 987, 987, 988, 988, 988, 988, 988, 988, 988, 988, 988, 988, 988, 988, 988, 988, 988, 989, 989, 989, 989, 989, 989, 989, 989, 989, 989, 989, 989, 989, 989, 989, 990, 990, 990, 990, 990, 990, 990, 990, 990, 990, 990, 990, 990, 990, 990, 990, 991, 991, 991, 991, 991, 991, 991, 991, 991, 991, 991, 991, 991, 991, 991, 991, 992, 992, 992, 992, 992, 992, 992, 992, 992, 992, 992, 992, 992, 992, 992, 992, 993, 993, 993, 993, 993, 993, 993, 993, 993, 993, 993, 993, 993, 993, 993, 993, 993, 994, 994, 994, 994, 994, 994, 994, 994, 994, 994, 994, 994, 994, 994, 994, 994, 994, 994, 995, 995, 995, 995, 995, 995, 995, 995, 995, 995, 995, 995, 995, 995, 995, 995, 995, 995, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 996, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 997, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 998, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 999, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1000, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1001, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1002, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1003, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1004, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1005, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1006, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1007, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1008, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1009, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1011, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1012, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1013, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1014, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1015, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1016, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1017, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1018, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1019, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1020, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1021, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1022, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023);
	
	signal int_x : integer range 0 to 4095;
	
    signal s_int_x, s_sat_x_conj, s_mux_x, s_sat_x: std_logic_vector(BitO-3 downto 0);
	signal lut_y, s_mux_a, s_mux_z : std_logic_vector(BitL downto 0);
	signal s_mux_z_ext : std_logic_vector(BitY-1 downto 0);
    signal sat_c, mux_c : std_logic;
	
	component N_MUX_2to1 is
		generic (Nbit : positive);
		port(	
			n_x : IN std_logic_vector;
			n_y : IN std_logic_vector;
			c : IN std_logic;
			n_z : OUT std_logic_vector
		);
	end component N_MUX_2to1;
	
	component N_DFF is
		generic (Nbit : positive);
		port (
			n_d : IN std_logic_vector;
			en : IN std_logic;
			clk : IN std_logic;
			resetn : IN std_logic;
			n_q : OUT std_logic_vector
		);
	end component N_DFF;
	
begin

	s_int_x <= x(BitO-3 downto 0);
    sat_c <= x(x'left) XOR x(x'left - 1); -- Control bit for first MUX
    mux_c <= x(x'left) AND x(x'left - 1); -- Control bit for second MUX
    
    -- Before LUT MUX for Saturation
	MUX_SAT : N_MUX_2to1
	generic map (Nbit => BitO-2)
	port map (
		n_x => s_int_x,
		n_y => x"FFF", -- 4095 in exadecimal
		c => sat_c,
		n_z => s_sat_x
	);
    
	s_sat_x_conj <= not(s_sat_x);
	
	-- Before LUT MUX for Optimization
	MUX_X : N_MUX_2to1
	generic map (Nbit => BitO-2)
	port map (
		n_x => s_sat_x,
		n_y => s_sat_x_conj,
		c => mux_c,
		n_z => s_mux_x
	);
		
	-- LUT index and value selected
	int_x <= to_integer(unsigned(s_mux_x));
	lut_y <= '1' & std_logic_vector(to_unsigned(SigmoidLUT(int_x), BitL));
	
	-- LUT Optimized MUX input A, subtracting lut_y to 1 (Rappresented by 1024)
	s_mux_a <= std_logic_vector(to_unsigned(2047, BitL+1) - unsigned(lut_y));
	
	-- After LUT MUX for Optimization
	MUX_Y : N_MUX_2to1
	generic map (Nbit => BitL+1)
	port map (
		n_x => lut_y,
		n_y => s_mux_a,
		c => x(x'left),
		n_z => s_mux_z
	);
	
	s_mux_z_ext <= (15 downto 11 => '0') & s_mux_z;
	
	DFF_Y : N_DFF
	generic map (Nbit => BitY)
	port map (
		n_d => s_mux_z_ext,
		en => '1',
		clk => clk,
		resetn => resetn,
		n_q => y
	);

end internal;